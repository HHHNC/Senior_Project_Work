version https://git-lfs.github.com/spec/v1
oid sha256:33e2dd63ebdf7756190d506c4eeba0559354f17585e6a9b1c06217fa14b14ad9
size 27018
